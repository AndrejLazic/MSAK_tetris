

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

ENTITY char_rom_def IS
  PORT (
    clka : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END char_rom_def;

ARCHITECTURE char_rom_def_a OF char_rom_def IS

  type t_char_rom  is array (0 to 2**9-1) of  std_logic_vector(7 downto 0);
  signal char_rom : t_char_rom := (
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00011000",
		"00111100",
		"01100110",
		"01111110",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01100000",
		"01100000",
		"01100110",
		"00111100",
		"00000000",
		"01111000",
		"01101100",
		"01100110",
		"01100110",
		"01100110",
		"01101100",
		"01111000",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111000",
		"01100000",
		"01100000",
		"01111110",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111000",
		"01100000",
		"01100000",
		"01100000",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01101110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01111110",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"00111100",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00111100",
		"00000000",
		"00011110",
		"00001100",
		"00001100",
		"00001100",
		"00001100",
		"01101100",
		"00111000",
		"00000000",
		"01100110",
		"01101100",
		"01111000",
		"01110000",
		"01111000",
		"01101100",
		"01100110",
		"00000000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01111110",
		"00000000",
		"01100011",
		"01110111",
		"01111111",
		"01101011",
		"01100011",
		"01100011",
		"01100011",
		"00000000",
		"01100110",
		"01110110",
		"01111110",
		"01111110",
		"01101110",
		"01100110",
		"01100110",
		"00000000",
		"00111100",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01100000",
		"01100000",
		"01100000",
		"00000000",
		"00111100",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00001110",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01111000",
		"01101100",
		"01100110",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"00111100",
		"00000110",
		"01100110",
		"00111100",
		"00000000",
		"01111110",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00000000",
		"01100011",
		"01100011",
		"01100011",
		"01101011",
		"01111111",
		"01110111",
		"01100011",
		"00000000",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00111100",
		"01100110",
		"01100110",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"01111110", --z start
		"00000110",
		"00001100",
		"00011000",
		"00110000",
		"01100000",
		"01111110",
		"00000000", --z end
		"00000000", -- kocka
		"00000000",
		"00111100",
		"00111100",
		"00111100",
		"00111100",
		"00000000",
		"00000000",-- kocka
		--ovde pocinju brojevi
		"00111100",
		"01100110",
		"01101110",
		"01110110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",--0
		"00011000",
		"00011000",
		"00111000",
		"00011000",
		"00011000",
		"00011000",
		"01111110",
		"00000000",--1
		"00111100",
		"01100110",
		"00000110",
		"00001100",
		"00110000",
		"01100000",
		"01111110",
		"00000000",--2
		"00111100",
		"01100110",
		"00000110",
		"00011100",
		"00000110",
		"01100110",
		"00111100",
		"00000000",--3
		"00000110",
		"00001110",
		"00011110",
		"01100110",
		"01111111",
		"00000110",
		"00000110",
		"00000000",--4
		"01111110",
		"01100000",
		"01111100",
		"00000110",
		"00000110",
		"01100110",
		"00111100",
		"00000000",--5
		"00111100",
		"01100110",
		"01100000",
		"01111100",
		"01100110",
		"01100110",
		"00111100",
		"00000000",--6
		"01111110",
		"01100110",
		"00001100",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",--7
		"00111100",
		"01100110",
		"01100110",
		"00111100",
		"01100110",
		"01100110",
		"00111100",
		"00000000",--8
		"00111100",
		"01100110",
		"00111110",
		"00111110",
		"00000110",
		"01100110",
		"00111100",  
		"00000000",--9
		others => "00000000"
	);
begin
	process (clka) begin
		if (rising_edge(clka)) then
			douta <= char_rom(conv_integer(addra));
		end if;
	end process;
  
END char_rom_def_a;
